module game_logic
#(
)
(
    input wire  enable,
    input wire  rst_n,

    input wire  plus_ten_score,

    output reg [13:0] score 
)






endmodule