module gw_gao(
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[13] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[12] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[11] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[10] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[9] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[8] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[7] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[6] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[5] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[4] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[3] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[2] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[1] ,
    \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[0] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[13] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[12] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[11] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[10] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[9] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[8] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[7] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[6] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[5] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[4] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[3] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[2] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[1] ,
    \lcd_data_wrap_inst/lcd_data_inst/high_score[0] ,
    \lcd_data_wrap_inst/game_over_finished ,
    lcd_clk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[13] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[12] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[11] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[10] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[9] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[8] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[7] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[6] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[5] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[4] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[3] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[2] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[1] ;
input \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[0] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[13] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[12] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[11] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[10] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[9] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[8] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[7] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[6] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[5] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[4] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[3] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[2] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[1] ;
input \lcd_data_wrap_inst/lcd_data_inst/high_score[0] ;
input \lcd_data_wrap_inst/game_over_finished ;
input lcd_clk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[13] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[12] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[11] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[10] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[9] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[8] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[7] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[6] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[5] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[4] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[3] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[2] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[1] ;
wire \lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[0] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[13] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[12] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[11] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[10] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[9] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[8] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[7] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[6] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[5] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[4] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[3] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[2] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[1] ;
wire \lcd_data_wrap_inst/lcd_data_inst/high_score[0] ;
wire \lcd_data_wrap_inst/game_over_finished ;
wire lcd_clk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i(\lcd_data_wrap_inst/game_over_finished ),
    .data_i({\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[13] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[12] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[11] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[10] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[9] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[8] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[7] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[6] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[5] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[4] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[3] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[2] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[1] ,\lcd_data_wrap_inst/lcd_data_inst/word_pixel_inst/score[0] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[13] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[12] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[11] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[10] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[9] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[8] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[7] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[6] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[5] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[4] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[3] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[2] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[1] ,\lcd_data_wrap_inst/lcd_data_inst/high_score[0] }),
    .clk_i(lcd_clk)
);

endmodule
